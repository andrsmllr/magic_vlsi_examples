magic
tech scmos
timestamp 1507236307
<< nwell >>
rect 0 0 24 16
<< ptransistor >>
rect 11 6 13 10
<< pdiffusion >>
rect 10 6 11 10
rect 13 6 14 10
<< pdcontact >>
rect 6 6 10 10
rect 14 6 18 10
<< polysilicon >>
rect 11 10 13 12
rect 11 0 13 6
<< polycontact >>
rect 13 0 17 4
<< metal1 >>
rect 3 6 6 10
rect 18 6 21 10
rect 14 4 17 6
<< labels >>
rlabel metal1 4 8 4 8 1 P
rlabel metal1 20 8 20 8 1 N
<< end >>
