* SPICE3 file created from transmissiongate.ext - technology: scmos

.option scale=0.25u

M1000 OUT CB IN Vdd pfet w=32 l=8
+  ad=640 pd=104 as=640 ps=104
M1001 OUT C IN GND nfet w=16 l=8
+  ad=320 pd=72 as=320 ps=72
C0 C GND 5.29fF
C1 CB Vdd 5.29fF
