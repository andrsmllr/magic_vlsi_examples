* SPICE3 file created from diode_nwpd.ext - technology: scmos

.option scale=0.05u

