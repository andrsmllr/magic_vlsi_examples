* SPICE3 file created from mux2.ext - technology: scmos

.option scale=0.05u

M1000 transmissiongate_0/OUT SB I0 Vdd pfet w=32 l=8
+  ad=640 pd=104 as=640 ps=104
M1001 transmissiongate_0/OUT S I0 GND nfet w=16 l=8
+  ad=320 pd=72 as=320 ps=72
M1002 transmissiongate_1/OUT S I1 Vdd pfet w=32 l=8
+  ad=640 pd=104 as=640 ps=104
M1003 transmissiongate_1/OUT SB I1 GND nfet w=16 l=8
+  ad=320 pd=72 as=320 ps=72
C0 Vdd 0 3.22fF
