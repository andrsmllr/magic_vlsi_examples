* SPICE3 file created from nor2.ext - technology: scmos

.option scale=0.25u

M1000 GND A OUT GND nfet w=16 l=12
+  ad=640 pd=144 as=640 ps=144
M1001 a_56_128# B Vdd Vdd pfet w=32 l=12
+  ad=1280 pd=208 as=640 ps=104
M1002 OUT B GND GND nfet w=16 l=12
+  ad=0 pd=0 as=0 ps=0
M1003 OUT A a_56_128# Vdd pfet w=32 l=12
+  ad=640 pd=104 as=0 ps=0
C0 Vdd A 7.95fF
C1 B GND 5.49fF
C2 A GND 4.09fF
C3 OUT GND 3.85fF
C4 B Vdd 2.94fF
