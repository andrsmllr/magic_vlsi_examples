magic
tech scmos
timestamp 1507279462
<< metal1 >>
rect -12 100 25 104
rect -12 78 0 82
rect -6 59 0 63
rect -12 52 25 56
rect -12 45 -4 49
rect -12 26 0 30
rect -12 11 -10 15
rect -6 11 0 15
rect -12 4 25 8
<< m2contact >>
rect -4 93 0 97
rect -10 59 -6 63
rect -4 45 0 49
rect -10 11 -6 15
<< metal2 >>
rect -10 15 -7 59
rect -3 49 0 93
use transmissiongate  transmissiongate_1
timestamp 1507277604
transform 1 0 0 0 -1 108
box 0 0 24 59
use transmissiongate  transmissiongate_0
timestamp 1507277604
transform 1 0 0 0 1 0
box 0 0 24 59
<< labels >>
rlabel metal1 -12 11 -11 15 3 S
rlabel metal1 -12 45 -11 49 3 SB
rlabel metal1 -12 26 -11 30 3 I0
rlabel metal1 -12 78 -11 82 3 I1
rlabel metal1 -2 102 -2 102 1 GND!
rlabel metal1 -5 54 -5 54 1 Vdd!
rlabel metal1 -3 6 -3 6 1 GND!
<< end >>
