magic
tech scmos
timestamp 1615325264
<< pwell >>
rect 0 0 43 26
<< nwell >>
rect 0 26 43 52
<< polysilicon >>
rect 11 40 14 42
rect 28 40 31 42
rect 11 24 14 32
rect 28 30 31 32
rect 21 27 31 30
rect 11 17 14 20
rect 28 17 31 27
rect 11 11 14 13
rect 28 11 31 13
<< ndiffusion >>
rect 10 13 11 17
rect 14 13 15 17
rect 27 13 28 17
rect 31 13 32 17
<< pdiffusion >>
rect 6 39 11 40
rect 10 33 11 39
rect 6 32 11 33
rect 14 39 19 40
rect 14 33 15 39
rect 14 32 19 33
rect 23 39 28 40
rect 27 33 28 39
rect 23 32 28 33
rect 31 39 36 40
rect 31 33 32 39
rect 31 32 36 33
<< metal1 >>
rect 0 44 4 48
rect 8 44 35 48
rect 39 44 43 48
rect 6 39 10 44
rect 19 33 23 39
rect 0 27 17 30
rect 33 26 36 33
rect 0 20 10 23
rect 24 23 43 26
rect 24 17 27 23
rect 19 13 23 17
rect 6 8 10 13
rect 32 8 36 13
rect 0 4 4 8
rect 8 4 35 8
rect 39 4 43 8
<< ntransistor >>
rect 11 13 14 17
rect 28 13 31 17
<< ptransistor >>
rect 11 32 14 40
rect 28 32 31 40
<< polycontact >>
rect 17 26 21 30
rect 10 20 14 24
<< ndcontact >>
rect 6 13 10 17
rect 15 13 19 17
rect 23 13 27 17
rect 32 13 36 17
<< pdcontact >>
rect 6 33 10 39
rect 15 33 19 39
rect 23 33 27 39
rect 32 33 36 39
<< psubstratepcontact >>
rect 4 4 8 8
rect 35 4 39 8
<< nsubstratencontact >>
rect 4 44 8 48
rect 35 44 39 48
<< labels >>
rlabel metal1 21 46 21 46 1 Vdd!
rlabel metal1 22 6 22 6 1 GND!
rlabel metal1 0 27 1 30 3 A
rlabel metal1 0 20 1 23 3 B
rlabel metal1 42 23 43 26 7 OUT
<< end >>
