magic
tech scmos
timestamp 1507281739
<< metal1 >>
rect -7 47 208 51
rect 205 34 208 38
rect -7 29 0 32
rect 49 29 53 32
rect -7 23 -4 26
rect 95 20 98 31
rect 148 29 150 32
rect 154 29 159 32
rect 148 28 152 29
rect 205 26 208 30
rect 156 20 159 26
rect -7 4 208 8
<< m2contact >>
rect 201 34 205 38
rect 42 28 46 32
rect -4 22 0 26
rect 49 22 53 26
rect 102 29 106 33
rect 150 29 154 33
rect 201 26 205 30
rect 102 22 106 26
rect 95 16 99 20
rect 155 16 159 20
<< metal2 >>
rect 150 34 201 38
rect 150 33 154 34
rect 46 29 102 32
rect 0 22 49 25
rect 106 23 205 26
rect 99 16 155 19
use nand2  nand2_0
timestamp 1507276308
transform 1 0 0 0 1 0
box 0 0 42 54
use nand2  nand2_1
timestamp 1507276308
transform 1 0 53 0 1 0
box 0 0 42 54
use nand2  nand2_2
timestamp 1507276308
transform 1 0 106 0 1 0
box 0 0 42 54
use nand2  nand2_3
timestamp 1507276308
transform 1 0 159 0 1 0
box 0 0 42 54
<< labels >>
rlabel metal1 -6 49 -6 49 3 Vdd!
rlabel metal1 -6 6 -6 6 3 GND!
rlabel metal1 -6 30 -6 30 3 D
rlabel metal1 -6 24 -6 24 3 E
rlabel metal1 207 34 208 38 7 Q
rlabel metal1 207 26 208 30 7 QB
<< end >>
