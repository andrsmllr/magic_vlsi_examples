magic
tech scmos
magscale 1 4
timestamp 1507277604
<< checkpaint >>
rect -104 232 197 233
rect -116 -8 212 232
<< nwell >>
rect 0 112 96 236
<< pwell >>
rect 0 0 96 112
<< ntransistor >>
rect 44 72 52 88
<< ptransistor >>
rect 44 136 52 168
<< ndiffusion >>
rect 40 72 44 88
rect 52 72 56 88
<< pdiffusion >>
rect 40 136 44 168
rect 52 136 56 168
<< ndcontact >>
rect 24 72 40 88
rect 56 72 72 88
<< pdcontact >>
rect 24 136 40 168
rect 56 136 72 168
<< psubstratepcontact >>
rect 16 16 32 32
rect 64 16 80 32
<< nsubstratencontact >>
rect 16 208 32 224
rect 64 208 80 224
<< polysilicon >>
rect 44 168 52 180
rect 44 128 52 136
rect 44 88 52 96
rect 44 60 52 72
<< polycontact >>
rect 40 180 56 196
rect 40 44 56 60
<< metal1 >>
rect 0 208 16 224
rect 32 208 64 224
rect 80 208 96 224
rect 0 180 40 196
rect 24 120 36 136
rect 0 104 36 120
rect 24 88 36 104
rect 60 120 72 136
rect 60 104 96 120
rect 60 88 72 104
rect 0 44 40 60
rect 0 16 16 32
rect 32 16 64 32
rect 80 16 96 32
<< labels >>
rlabel metal1 48 24 48 24 1 GND!
rlabel metal1 8 52 8 52 1 C
rlabel metal1 8 188 8 188 1 CB
rlabel metal1 44 216 44 216 1 Vdd!
rlabel metal1 0 104 4 120 3 IN
rlabel metal1 92 104 96 120 7 OUT
<< end >>
