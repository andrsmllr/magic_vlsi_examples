magic
tech scmos
timestamp 1507235735
<< pwell >>
rect 0 0 25 17
<< ntransistor >>
rect 11 6 14 11
<< ndiffusion >>
rect 10 6 11 11
rect 14 6 15 11
<< ndcontact >>
rect 6 6 10 11
rect 15 6 19 11
<< polysilicon >>
rect 11 11 14 17
rect 11 4 14 6
<< polycontact >>
rect 7 13 11 17
<< metal1 >>
rect 7 11 10 13
rect 3 7 6 10
rect 19 7 22 10
<< labels >>
rlabel metal1 4 8 4 8 3 P
rlabel metal1 20 8 20 8 1 N
<< end >>
